package types;

typedef logic[31:0] u32; 
typedef logic[15:0] u16;
typedef logic[ 7:0] u8;
typedef logic[ 3:0] u4;   







endpackage